VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_scoreboard
  CLASS BLOCK ;
  FOREIGN user_proj_scoreboard ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 3000.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2831.560 4.000 2832.160 ;
    END
  END io_in[0]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2498.360 4.000 2498.960 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2165.160 4.000 2165.760 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1831.960 4.000 1832.560 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1498.760 4.000 1499.360 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 1165.560 4.000 1166.160 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 832.360 4.000 832.960 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.160 4.000 499.760 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END io_in[8]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 2876.440 200.000 2877.040 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 1652.440 200.000 1653.040 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 1530.040 200.000 1530.640 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 1407.640 200.000 1408.240 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 1285.240 200.000 1285.840 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 1162.840 200.000 1163.440 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 1040.440 200.000 1041.040 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 918.040 200.000 918.640 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 795.640 200.000 796.240 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 673.240 200.000 673.840 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 550.840 200.000 551.440 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 2754.040 200.000 2754.640 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 428.440 200.000 429.040 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 306.040 200.000 306.640 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 183.640 200.000 184.240 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 61.240 200.000 61.840 ;
    END
  END io_oeb[23]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 2631.640 200.000 2632.240 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 2509.240 200.000 2509.840 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 2386.840 200.000 2387.440 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 2264.440 200.000 2265.040 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 2142.040 200.000 2142.640 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 2019.640 200.000 2020.240 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 1897.240 200.000 1897.840 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 1774.840 200.000 1775.440 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 2937.640 200.000 2938.240 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 1713.640 200.000 1714.240 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 1591.240 200.000 1591.840 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 1468.840 200.000 1469.440 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 1346.440 200.000 1347.040 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 1224.040 200.000 1224.640 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 1101.640 200.000 1102.240 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 979.240 200.000 979.840 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 856.840 200.000 857.440 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 734.440 200.000 735.040 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 612.040 200.000 612.640 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 2815.240 200.000 2815.840 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 489.640 200.000 490.240 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 367.240 200.000 367.840 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 244.840 200.000 245.440 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 122.440 200.000 123.040 ;
    END
  END io_out[23]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 2692.840 200.000 2693.440 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 2570.440 200.000 2571.040 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 2448.040 200.000 2448.640 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 2325.640 200.000 2326.240 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 2203.240 200.000 2203.840 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 2080.840 200.000 2081.440 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 1958.440 200.000 1959.040 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 196.000 1836.040 200.000 1836.640 ;
    END
  END io_out[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 2986.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 2986.800 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 2986.800 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.869400 ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 149.590 0.000 149.870 4.000 ;
    END
  END wb_rst_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.120 2986.645 ;
      LAYER met1 ;
        RECT 4.670 10.640 196.350 2986.800 ;
      LAYER met2 ;
        RECT 4.690 4.280 196.320 2986.745 ;
        RECT 4.690 4.000 49.490 4.280 ;
        RECT 50.330 4.000 149.310 4.280 ;
        RECT 150.150 4.000 196.320 4.280 ;
      LAYER met3 ;
        RECT 4.000 2938.640 196.000 2986.725 ;
        RECT 4.000 2937.240 195.600 2938.640 ;
        RECT 4.000 2877.440 196.000 2937.240 ;
        RECT 4.000 2876.040 195.600 2877.440 ;
        RECT 4.000 2832.560 196.000 2876.040 ;
        RECT 4.400 2831.160 196.000 2832.560 ;
        RECT 4.000 2816.240 196.000 2831.160 ;
        RECT 4.000 2814.840 195.600 2816.240 ;
        RECT 4.000 2755.040 196.000 2814.840 ;
        RECT 4.000 2753.640 195.600 2755.040 ;
        RECT 4.000 2693.840 196.000 2753.640 ;
        RECT 4.000 2692.440 195.600 2693.840 ;
        RECT 4.000 2632.640 196.000 2692.440 ;
        RECT 4.000 2631.240 195.600 2632.640 ;
        RECT 4.000 2571.440 196.000 2631.240 ;
        RECT 4.000 2570.040 195.600 2571.440 ;
        RECT 4.000 2510.240 196.000 2570.040 ;
        RECT 4.000 2508.840 195.600 2510.240 ;
        RECT 4.000 2499.360 196.000 2508.840 ;
        RECT 4.400 2497.960 196.000 2499.360 ;
        RECT 4.000 2449.040 196.000 2497.960 ;
        RECT 4.000 2447.640 195.600 2449.040 ;
        RECT 4.000 2387.840 196.000 2447.640 ;
        RECT 4.000 2386.440 195.600 2387.840 ;
        RECT 4.000 2326.640 196.000 2386.440 ;
        RECT 4.000 2325.240 195.600 2326.640 ;
        RECT 4.000 2265.440 196.000 2325.240 ;
        RECT 4.000 2264.040 195.600 2265.440 ;
        RECT 4.000 2204.240 196.000 2264.040 ;
        RECT 4.000 2202.840 195.600 2204.240 ;
        RECT 4.000 2166.160 196.000 2202.840 ;
        RECT 4.400 2164.760 196.000 2166.160 ;
        RECT 4.000 2143.040 196.000 2164.760 ;
        RECT 4.000 2141.640 195.600 2143.040 ;
        RECT 4.000 2081.840 196.000 2141.640 ;
        RECT 4.000 2080.440 195.600 2081.840 ;
        RECT 4.000 2020.640 196.000 2080.440 ;
        RECT 4.000 2019.240 195.600 2020.640 ;
        RECT 4.000 1959.440 196.000 2019.240 ;
        RECT 4.000 1958.040 195.600 1959.440 ;
        RECT 4.000 1898.240 196.000 1958.040 ;
        RECT 4.000 1896.840 195.600 1898.240 ;
        RECT 4.000 1837.040 196.000 1896.840 ;
        RECT 4.000 1835.640 195.600 1837.040 ;
        RECT 4.000 1832.960 196.000 1835.640 ;
        RECT 4.400 1831.560 196.000 1832.960 ;
        RECT 4.000 1775.840 196.000 1831.560 ;
        RECT 4.000 1774.440 195.600 1775.840 ;
        RECT 4.000 1714.640 196.000 1774.440 ;
        RECT 4.000 1713.240 195.600 1714.640 ;
        RECT 4.000 1653.440 196.000 1713.240 ;
        RECT 4.000 1652.040 195.600 1653.440 ;
        RECT 4.000 1592.240 196.000 1652.040 ;
        RECT 4.000 1590.840 195.600 1592.240 ;
        RECT 4.000 1531.040 196.000 1590.840 ;
        RECT 4.000 1529.640 195.600 1531.040 ;
        RECT 4.000 1499.760 196.000 1529.640 ;
        RECT 4.400 1498.360 196.000 1499.760 ;
        RECT 4.000 1469.840 196.000 1498.360 ;
        RECT 4.000 1468.440 195.600 1469.840 ;
        RECT 4.000 1408.640 196.000 1468.440 ;
        RECT 4.000 1407.240 195.600 1408.640 ;
        RECT 4.000 1347.440 196.000 1407.240 ;
        RECT 4.000 1346.040 195.600 1347.440 ;
        RECT 4.000 1286.240 196.000 1346.040 ;
        RECT 4.000 1284.840 195.600 1286.240 ;
        RECT 4.000 1225.040 196.000 1284.840 ;
        RECT 4.000 1223.640 195.600 1225.040 ;
        RECT 4.000 1166.560 196.000 1223.640 ;
        RECT 4.400 1165.160 196.000 1166.560 ;
        RECT 4.000 1163.840 196.000 1165.160 ;
        RECT 4.000 1162.440 195.600 1163.840 ;
        RECT 4.000 1102.640 196.000 1162.440 ;
        RECT 4.000 1101.240 195.600 1102.640 ;
        RECT 4.000 1041.440 196.000 1101.240 ;
        RECT 4.000 1040.040 195.600 1041.440 ;
        RECT 4.000 980.240 196.000 1040.040 ;
        RECT 4.000 978.840 195.600 980.240 ;
        RECT 4.000 919.040 196.000 978.840 ;
        RECT 4.000 917.640 195.600 919.040 ;
        RECT 4.000 857.840 196.000 917.640 ;
        RECT 4.000 856.440 195.600 857.840 ;
        RECT 4.000 833.360 196.000 856.440 ;
        RECT 4.400 831.960 196.000 833.360 ;
        RECT 4.000 796.640 196.000 831.960 ;
        RECT 4.000 795.240 195.600 796.640 ;
        RECT 4.000 735.440 196.000 795.240 ;
        RECT 4.000 734.040 195.600 735.440 ;
        RECT 4.000 674.240 196.000 734.040 ;
        RECT 4.000 672.840 195.600 674.240 ;
        RECT 4.000 613.040 196.000 672.840 ;
        RECT 4.000 611.640 195.600 613.040 ;
        RECT 4.000 551.840 196.000 611.640 ;
        RECT 4.000 550.440 195.600 551.840 ;
        RECT 4.000 500.160 196.000 550.440 ;
        RECT 4.400 498.760 196.000 500.160 ;
        RECT 4.000 490.640 196.000 498.760 ;
        RECT 4.000 489.240 195.600 490.640 ;
        RECT 4.000 429.440 196.000 489.240 ;
        RECT 4.000 428.040 195.600 429.440 ;
        RECT 4.000 368.240 196.000 428.040 ;
        RECT 4.000 366.840 195.600 368.240 ;
        RECT 4.000 307.040 196.000 366.840 ;
        RECT 4.000 305.640 195.600 307.040 ;
        RECT 4.000 245.840 196.000 305.640 ;
        RECT 4.000 244.440 195.600 245.840 ;
        RECT 4.000 184.640 196.000 244.440 ;
        RECT 4.000 183.240 195.600 184.640 ;
        RECT 4.000 166.960 196.000 183.240 ;
        RECT 4.400 165.560 196.000 166.960 ;
        RECT 4.000 123.440 196.000 165.560 ;
        RECT 4.000 122.040 195.600 123.440 ;
        RECT 4.000 62.240 196.000 122.040 ;
        RECT 4.000 60.840 195.600 62.240 ;
        RECT 4.000 10.715 196.000 60.840 ;
      LAYER met4 ;
        RECT 113.455 17.175 174.240 1711.385 ;
        RECT 176.640 17.175 185.545 1711.385 ;
  END
END user_proj_scoreboard
END LIBRARY

