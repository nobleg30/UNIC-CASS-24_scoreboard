magic
tech sky130A
magscale 1 2
timestamp 1729621189
<< obsli1 >>
rect 1104 2159 38824 597329
<< obsm1 >>
rect 934 2128 39270 597360
<< metal2 >>
rect 9954 0 10010 800
rect 29918 0 29974 800
<< obsm2 >>
rect 938 856 39264 597349
rect 938 800 9898 856
rect 10066 800 29862 856
rect 30030 800 39264 856
<< metal3 >>
rect 39200 587528 40000 587648
rect 39200 575288 40000 575408
rect 0 566312 800 566432
rect 39200 563048 40000 563168
rect 39200 550808 40000 550928
rect 39200 538568 40000 538688
rect 39200 526328 40000 526448
rect 39200 514088 40000 514208
rect 39200 501848 40000 501968
rect 0 499672 800 499792
rect 39200 489608 40000 489728
rect 39200 477368 40000 477488
rect 39200 465128 40000 465248
rect 39200 452888 40000 453008
rect 39200 440648 40000 440768
rect 0 433032 800 433152
rect 39200 428408 40000 428528
rect 39200 416168 40000 416288
rect 39200 403928 40000 404048
rect 39200 391688 40000 391808
rect 39200 379448 40000 379568
rect 39200 367208 40000 367328
rect 0 366392 800 366512
rect 39200 354968 40000 355088
rect 39200 342728 40000 342848
rect 39200 330488 40000 330608
rect 39200 318248 40000 318368
rect 39200 306008 40000 306128
rect 0 299752 800 299872
rect 39200 293768 40000 293888
rect 39200 281528 40000 281648
rect 39200 269288 40000 269408
rect 39200 257048 40000 257168
rect 39200 244808 40000 244928
rect 0 233112 800 233232
rect 39200 232568 40000 232688
rect 39200 220328 40000 220448
rect 39200 208088 40000 208208
rect 39200 195848 40000 195968
rect 39200 183608 40000 183728
rect 39200 171368 40000 171488
rect 0 166472 800 166592
rect 39200 159128 40000 159248
rect 39200 146888 40000 147008
rect 39200 134648 40000 134768
rect 39200 122408 40000 122528
rect 39200 110168 40000 110288
rect 0 99832 800 99952
rect 39200 97928 40000 98048
rect 39200 85688 40000 85808
rect 39200 73448 40000 73568
rect 39200 61208 40000 61328
rect 39200 48968 40000 49088
rect 39200 36728 40000 36848
rect 0 33192 800 33312
rect 39200 24488 40000 24608
rect 39200 12248 40000 12368
<< obsm3 >>
rect 800 587728 39200 597345
rect 800 587448 39120 587728
rect 800 575488 39200 587448
rect 800 575208 39120 575488
rect 800 566512 39200 575208
rect 880 566232 39200 566512
rect 800 563248 39200 566232
rect 800 562968 39120 563248
rect 800 551008 39200 562968
rect 800 550728 39120 551008
rect 800 538768 39200 550728
rect 800 538488 39120 538768
rect 800 526528 39200 538488
rect 800 526248 39120 526528
rect 800 514288 39200 526248
rect 800 514008 39120 514288
rect 800 502048 39200 514008
rect 800 501768 39120 502048
rect 800 499872 39200 501768
rect 880 499592 39200 499872
rect 800 489808 39200 499592
rect 800 489528 39120 489808
rect 800 477568 39200 489528
rect 800 477288 39120 477568
rect 800 465328 39200 477288
rect 800 465048 39120 465328
rect 800 453088 39200 465048
rect 800 452808 39120 453088
rect 800 440848 39200 452808
rect 800 440568 39120 440848
rect 800 433232 39200 440568
rect 880 432952 39200 433232
rect 800 428608 39200 432952
rect 800 428328 39120 428608
rect 800 416368 39200 428328
rect 800 416088 39120 416368
rect 800 404128 39200 416088
rect 800 403848 39120 404128
rect 800 391888 39200 403848
rect 800 391608 39120 391888
rect 800 379648 39200 391608
rect 800 379368 39120 379648
rect 800 367408 39200 379368
rect 800 367128 39120 367408
rect 800 366592 39200 367128
rect 880 366312 39200 366592
rect 800 355168 39200 366312
rect 800 354888 39120 355168
rect 800 342928 39200 354888
rect 800 342648 39120 342928
rect 800 330688 39200 342648
rect 800 330408 39120 330688
rect 800 318448 39200 330408
rect 800 318168 39120 318448
rect 800 306208 39200 318168
rect 800 305928 39120 306208
rect 800 299952 39200 305928
rect 880 299672 39200 299952
rect 800 293968 39200 299672
rect 800 293688 39120 293968
rect 800 281728 39200 293688
rect 800 281448 39120 281728
rect 800 269488 39200 281448
rect 800 269208 39120 269488
rect 800 257248 39200 269208
rect 800 256968 39120 257248
rect 800 245008 39200 256968
rect 800 244728 39120 245008
rect 800 233312 39200 244728
rect 880 233032 39200 233312
rect 800 232768 39200 233032
rect 800 232488 39120 232768
rect 800 220528 39200 232488
rect 800 220248 39120 220528
rect 800 208288 39200 220248
rect 800 208008 39120 208288
rect 800 196048 39200 208008
rect 800 195768 39120 196048
rect 800 183808 39200 195768
rect 800 183528 39120 183808
rect 800 171568 39200 183528
rect 800 171288 39120 171568
rect 800 166672 39200 171288
rect 880 166392 39200 166672
rect 800 159328 39200 166392
rect 800 159048 39120 159328
rect 800 147088 39200 159048
rect 800 146808 39120 147088
rect 800 134848 39200 146808
rect 800 134568 39120 134848
rect 800 122608 39200 134568
rect 800 122328 39120 122608
rect 800 110368 39200 122328
rect 800 110088 39120 110368
rect 800 100032 39200 110088
rect 880 99752 39200 100032
rect 800 98128 39200 99752
rect 800 97848 39120 98128
rect 800 85888 39200 97848
rect 800 85608 39120 85888
rect 800 73648 39200 85608
rect 800 73368 39120 73648
rect 800 61408 39200 73368
rect 800 61128 39120 61408
rect 800 49168 39200 61128
rect 800 48888 39120 49168
rect 800 36928 39200 48888
rect 800 36648 39120 36928
rect 800 33392 39200 36648
rect 880 33112 39200 33392
rect 800 24688 39200 33112
rect 800 24408 39120 24688
rect 800 12448 39200 24408
rect 800 12168 39120 12448
rect 800 2143 39200 12168
<< metal4 >>
rect 4208 2128 4528 597360
rect 19568 2128 19888 597360
rect 34928 2128 35248 597360
<< obsm4 >>
rect 22691 3435 34848 342277
rect 35328 3435 37109 342277
<< labels >>
rlabel metal3 s 0 566312 800 566432 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 0 499672 800 499792 6 io_in[1]
port 2 nsew signal input
rlabel metal3 s 0 433032 800 433152 6 io_in[2]
port 3 nsew signal input
rlabel metal3 s 0 366392 800 366512 6 io_in[3]
port 4 nsew signal input
rlabel metal3 s 0 299752 800 299872 6 io_in[4]
port 5 nsew signal input
rlabel metal3 s 0 233112 800 233232 6 io_in[5]
port 6 nsew signal input
rlabel metal3 s 0 166472 800 166592 6 io_in[6]
port 7 nsew signal input
rlabel metal3 s 0 99832 800 99952 6 io_in[7]
port 8 nsew signal input
rlabel metal3 s 0 33192 800 33312 6 io_in[8]
port 9 nsew signal input
rlabel metal3 s 39200 575288 40000 575408 6 io_oeb[0]
port 10 nsew signal output
rlabel metal3 s 39200 330488 40000 330608 6 io_oeb[10]
port 11 nsew signal output
rlabel metal3 s 39200 306008 40000 306128 6 io_oeb[11]
port 12 nsew signal output
rlabel metal3 s 39200 281528 40000 281648 6 io_oeb[12]
port 13 nsew signal output
rlabel metal3 s 39200 257048 40000 257168 6 io_oeb[13]
port 14 nsew signal output
rlabel metal3 s 39200 232568 40000 232688 6 io_oeb[14]
port 15 nsew signal output
rlabel metal3 s 39200 208088 40000 208208 6 io_oeb[15]
port 16 nsew signal output
rlabel metal3 s 39200 183608 40000 183728 6 io_oeb[16]
port 17 nsew signal output
rlabel metal3 s 39200 159128 40000 159248 6 io_oeb[17]
port 18 nsew signal output
rlabel metal3 s 39200 134648 40000 134768 6 io_oeb[18]
port 19 nsew signal output
rlabel metal3 s 39200 110168 40000 110288 6 io_oeb[19]
port 20 nsew signal output
rlabel metal3 s 39200 550808 40000 550928 6 io_oeb[1]
port 21 nsew signal output
rlabel metal3 s 39200 85688 40000 85808 6 io_oeb[20]
port 22 nsew signal output
rlabel metal3 s 39200 61208 40000 61328 6 io_oeb[21]
port 23 nsew signal output
rlabel metal3 s 39200 36728 40000 36848 6 io_oeb[22]
port 24 nsew signal output
rlabel metal3 s 39200 12248 40000 12368 6 io_oeb[23]
port 25 nsew signal output
rlabel metal3 s 39200 526328 40000 526448 6 io_oeb[2]
port 26 nsew signal output
rlabel metal3 s 39200 501848 40000 501968 6 io_oeb[3]
port 27 nsew signal output
rlabel metal3 s 39200 477368 40000 477488 6 io_oeb[4]
port 28 nsew signal output
rlabel metal3 s 39200 452888 40000 453008 6 io_oeb[5]
port 29 nsew signal output
rlabel metal3 s 39200 428408 40000 428528 6 io_oeb[6]
port 30 nsew signal output
rlabel metal3 s 39200 403928 40000 404048 6 io_oeb[7]
port 31 nsew signal output
rlabel metal3 s 39200 379448 40000 379568 6 io_oeb[8]
port 32 nsew signal output
rlabel metal3 s 39200 354968 40000 355088 6 io_oeb[9]
port 33 nsew signal output
rlabel metal3 s 39200 587528 40000 587648 6 io_out[0]
port 34 nsew signal output
rlabel metal3 s 39200 342728 40000 342848 6 io_out[10]
port 35 nsew signal output
rlabel metal3 s 39200 318248 40000 318368 6 io_out[11]
port 36 nsew signal output
rlabel metal3 s 39200 293768 40000 293888 6 io_out[12]
port 37 nsew signal output
rlabel metal3 s 39200 269288 40000 269408 6 io_out[13]
port 38 nsew signal output
rlabel metal3 s 39200 244808 40000 244928 6 io_out[14]
port 39 nsew signal output
rlabel metal3 s 39200 220328 40000 220448 6 io_out[15]
port 40 nsew signal output
rlabel metal3 s 39200 195848 40000 195968 6 io_out[16]
port 41 nsew signal output
rlabel metal3 s 39200 171368 40000 171488 6 io_out[17]
port 42 nsew signal output
rlabel metal3 s 39200 146888 40000 147008 6 io_out[18]
port 43 nsew signal output
rlabel metal3 s 39200 122408 40000 122528 6 io_out[19]
port 44 nsew signal output
rlabel metal3 s 39200 563048 40000 563168 6 io_out[1]
port 45 nsew signal output
rlabel metal3 s 39200 97928 40000 98048 6 io_out[20]
port 46 nsew signal output
rlabel metal3 s 39200 73448 40000 73568 6 io_out[21]
port 47 nsew signal output
rlabel metal3 s 39200 48968 40000 49088 6 io_out[22]
port 48 nsew signal output
rlabel metal3 s 39200 24488 40000 24608 6 io_out[23]
port 49 nsew signal output
rlabel metal3 s 39200 538568 40000 538688 6 io_out[2]
port 50 nsew signal output
rlabel metal3 s 39200 514088 40000 514208 6 io_out[3]
port 51 nsew signal output
rlabel metal3 s 39200 489608 40000 489728 6 io_out[4]
port 52 nsew signal output
rlabel metal3 s 39200 465128 40000 465248 6 io_out[5]
port 53 nsew signal output
rlabel metal3 s 39200 440648 40000 440768 6 io_out[6]
port 54 nsew signal output
rlabel metal3 s 39200 416168 40000 416288 6 io_out[7]
port 55 nsew signal output
rlabel metal3 s 39200 391688 40000 391808 6 io_out[8]
port 56 nsew signal output
rlabel metal3 s 39200 367208 40000 367328 6 io_out[9]
port 57 nsew signal output
rlabel metal4 s 4208 2128 4528 597360 6 vccd1
port 58 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 597360 6 vccd1
port 58 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 597360 6 vssd1
port 59 nsew ground bidirectional
rlabel metal2 s 9954 0 10010 800 6 wb_clk_i
port 60 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 wb_rst_i
port 61 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 40000 600000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 18398158
string GDS_FILE /home/ngk/unic_cass_ic/uniccass_example/openlane/user_proj_scoreboard/runs/24_10_22_23_46/results/signoff/user_proj_scoreboard.magic.gds
string GDS_START 1015506
<< end >>

